package configure;

	parameter start_addr = 32'h0;

	parameter memory_depth = 12;

endpackage
