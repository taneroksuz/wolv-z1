timeunit 1ns;
timeprecision 1ps;

module test_cpu
(
	input reset,
	input clock
);

endmodule
