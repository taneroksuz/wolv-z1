module fetch_stage();

endmodule
