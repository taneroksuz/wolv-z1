import wires::*;
import functions::*;

module bit_clmul
(
  input logic rst,
  input logic clk,
  input bit_clmul_in_type bit_clmul_in,
  output bit_clmul_out_type bit_clmul_out
);
  timeunit 1ns;
  timeprecision 1ps;

  always_comb begin


  end

endmodule
