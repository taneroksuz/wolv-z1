module decode_stage();

endmodule
