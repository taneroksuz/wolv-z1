module wires();

endmodule
